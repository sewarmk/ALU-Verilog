module checkgreater(g,A,B);
input [7:0]A;
input [7:0]B;
wire [7:0]o;
wire [7:0]w;
wire [7:0]p;
wire [7:0]i;
wire [7:0]v;
wire j;
output g;
onescomplement ones500(o,B);
and a1(w[0],A[7],o[7]);
and a2(w[1],A[6],o[6]);
and a3(w[2],A[5],o[5]);
and a4(w[3],A[4],o[4]);
and a5(w[4],A[3],o[3]);
and a6(w[5],A[2],o[2]);
and a7(w[6],A[1],o[1]);
and a8(w[7],A[0],o[0]);
xnor x1(p[0],A[7],B[7]);
xnor x2(p[1],A[6],B[6]);
xnor x3(p[2],A[5],B[5]);
xnor x4(p[3],A[4],B[4]);
xnor x5(p[4],A[3],B[3]);
xnor x6(p[5],A[2],B[2]);
xnor x7(p[6],A[1],B[1]);
xnor x8(p[7],A[0],B[0]);
assign v[0]=w[0];
and t1(v[1],p[0],w[1]);
and t2(v[2],p[0],p[1],w[2]);
and t3(v[3],p[0],p[1],p[2],w[3]);
and t5(v[4],p[0],p[1],p[2],p[3],w[4]);
and t6(v[5],p[0],p[1],p[2],p[3],p[4],w[5]);
and t7(v[6],p[0],p[1],p[2],p[3],p[4],p[5],w[6]);
and t8(v[7],p[0],p[1],p[2],p[3],p[4],p[5],p[6],w[7]);

or q1(j,v[0],v[1],v[2],v[3],v[4],v[5],v[6],v[7]);
assign g = (j)?1'b1:1'b0;
endmodule 